----------------------------------------------------------------------------------
-- Company: UC3M
-- Engineer: Alejandro Estaire Martin
-- 
-- Create Date: 27.05.2025 20:15:37
-- Design Name: 
-- Module Name: gen_seno - Behavioral
-- Project Name: Audiometry
-- Target Devices: Basys3 & Pmod I2S2
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity gen_seno is
  port(
    clk          : in  std_logic;
    tick         : in  std_logic;
    new_freq     : in  std_logic;
    cuenta_max   : in  unsigned(14 downto 0);
    gen_seno_out : out std_logic_vector(23 downto 0)
  );
end gen_seno;

architecture Behavioral of gen_seno is
  type seno_lut_type is array(0 to 4095) of signed(23 downto 0);
  signal seno_lut : seno_lut_type := (
    -- Cargar desde archivo externo generado en Python
    x"000000", x"003243", x"006487", x"0096CB", x"00C90F", x"00FB53", x"012D96", x"015FDA", x"01921D", x"01C45F",
x"01F6A2", x"0228E4", x"025B26", x"028D68", x"02BFA9", x"02F1EA", x"03242A", x"03566A", x"0388A9", x"03BAE8",
x"03ED26", x"041F64", x"0451A1", x"0483DD", x"04B619", x"04E854", x"051A8E", x"054CC7", x"057F00", x"05B137",
x"05E36E", x"0615A4", x"0647D9", x"067A0D", x"06AC40", x"06DE72", x"0710A3", x"0742D3", x"077501", x"07A72F",
x"07D95B", x"080B86", x"083DB0", x"086FD9", x"08A200", x"08D426", x"09064B", x"09386E", x"096A90", x"099CB0",
x"09CECF", x"0A00EC", x"0A3308", x"0A6522", x"0A973B", x"0AC952", x"0AFB67", x"0B2D7B", x"0B5F8D", x"0B919D",
x"0BC3AC", x"0BF5B8", x"0C27C3", x"0C59CC", x"0C8BD3", x"0CBDD8", x"0CEFDB", x"0D21DC", x"0D53DB", x"0D85D8",
x"0DB7D3", x"0DE9CC", x"0E1BC2", x"0E4DB7", x"0E7FA9", x"0EB199", x"0EE387", x"0F1572", x"0F475B", x"0F7942",
x"0FAB27", x"0FDD09", x"100EE8", x"1040C5", x"1072A0", x"10A478", x"10D64D", x"110820", x"1139F0", x"116BBE",
x"119D89", x"11CF51", x"120116", x"1232D9", x"126499", x"129656", x"12C810", x"12F9C7", x"132B7B", x"135D2D",
x"138EDB", x"13C086", x"13F22F", x"1423D4", x"145576", x"148715", x"14B8B1", x"14EA49", x"151BDF", x"154D71",
x"157F00", x"15B08B", x"15E214", x"161398", x"16451A", x"167698", x"16A812", x"16D989", x"170AFD", x"173C6D",
x"176DD9", x"179F42", x"17D0A7", x"180208", x"183366", x"1864C0", x"189616", x"18C769", x"18F8B8", x"192A02",
x"195B49", x"198C8C", x"19BDCB", x"19EF06", x"1A203D", x"1A5170", x"1A829F", x"1AB3CA", x"1AE4F1", x"1B1614",
x"1B4732", x"1B784C", x"1BA962", x"1BDA74", x"1C0B82", x"1C3C8B", x"1C6D90", x"1C9E90", x"1CCF8C", x"1D0084",
x"1D3177", x"1D6265", x"1D934F", x"1DC435", x"1DF516", x"1E25F2", x"1E56C9", x"1E879C", x"1EB86B", x"1EE934",
x"1F19F9", x"1F4AB9", x"1F7B74", x"1FAC2A", x"1FDCDB", x"200D88", x"203E2F", x"206ED2", x"209F6F", x"20D008",
x"21009B", x"21312A", x"2161B3", x"219237", x"21C2B6", x"21F330", x"2223A4", x"225413", x"22847D", x"22B4E2",
x"22E541", x"23159B", x"2345EF", x"23763E", x"23A688", x"23D6CC", x"24070A", x"243743", x"246777", x"2497A4",
x"24C7CC", x"24F7EF", x"25280C", x"255823", x"258834", x"25B83F", x"25E845", x"261845", x"26483F", x"267833",
x"26A821", x"26D809", x"2707EB", x"2737C7", x"27679D", x"27976D", x"27C737", x"27F6FB", x"2826B8", x"285670",
x"288621", x"28B5CC", x"28E570", x"29150F", x"2944A7", x"297438", x"29A3C4", x"29D349", x"2A02C7", x"2A323F",
x"2A61B0", x"2A911B", x"2AC07F", x"2AEFDD", x"2B1F34", x"2B4E85", x"2B7DCE", x"2BAD11", x"2BDC4E", x"2C0B83",
x"2C3AB2", x"2C69DA", x"2C98FB", x"2CC815", x"2CF728", x"2D2635", x"2D553A", x"2D8439", x"2DB330", x"2DE220",
x"2E110A", x"2E3FEC", x"2E6EC7", x"2E9D9B", x"2ECC67", x"2EFB2D", x"2F29EB", x"2F58A2", x"2F8752", x"2FB5FA",
x"2FE49B", x"301334", x"3041C7", x"307051", x"309ED4", x"30CD50", x"30FBC4", x"312A31", x"315896", x"3186F4",
x"31B549", x"31E398", x"3211DE", x"32401D", x"326E54", x"329C83", x"32CAAB", x"32F8CA", x"3326E2", x"3354F2",
x"3382FA", x"33B0FA", x"33DEF2", x"340CE2", x"343ACA", x"3468AA", x"349681", x"34C451", x"34F219", x"351FD8",
x"354D8F", x"357B3E", x"35A8E5", x"35D684", x"36041A", x"3631A8", x"365F2D", x"368CAA", x"36BA1F", x"36E78B",
x"3714EF", x"37424B", x"376F9D", x"379CE8", x"37CA29", x"37F762", x"382493", x"3851BB", x"387EDA", x"38ABF0",
x"38D8FE", x"390603", x"3932FF", x"395FF2", x"398CDC", x"39B9BE", x"39E696", x"3A1366", x"3A402D", x"3A6CEB",
x"3A999F", x"3AC64B", x"3AF2EE", x"3B1F87", x"3B4C18", x"3B789F", x"3BA51D", x"3BD192", x"3BFDFE", x"3C2A60",
x"3C56B9", x"3C8309", x"3CAF50", x"3CDB8D", x"3D07C1", x"3D33EB", x"3D600C", x"3D8C24", x"3DB832", x"3DE436",
x"3E1031", x"3E3C22", x"3E680A", x"3E93E8", x"3EBFBD", x"3EEB88", x"3F1749", x"3F4300", x"3F6EAE", x"3F9A52",
x"3FC5EC", x"3FF17C", x"401D02", x"40487F", x"4073F1", x"409F5A", x"40CAB8", x"40F60D", x"412158", x"414C98",
x"4177CF", x"41A2FB", x"41CE1D", x"41F936", x"422443", x"424F47", x"427A41", x"42A530", x"42D015", x"42FAF0",
x"4325C0", x"435086", x"437B42", x"43A5F3", x"43D09A", x"43FB36", x"4425C8", x"44504F", x"447ACC", x"44A53F",
x"44CFA6", x"44FA03", x"452456", x"454E9D", x"4578DB", x"45A30D", x"45CD35", x"45F751", x"462163", x"464B6B",
x"467567", x"469F59", x"46C93F", x"46F31B", x"471CEC", x"4746B2", x"47706D", x"479A1C", x"47C3C1", x"47ED5B",
x"4816E9", x"48406D", x"4869E5", x"489353", x"48BCB5", x"48E60B", x"490F57", x"493897", x"4961CC", x"498AF6",
x"49B414", x"49DD27", x"4A062F", x"4A2F2B", x"4A581C", x"4A8101", x"4AA9DB", x"4AD2A9", x"4AFB6C", x"4B2423",
x"4B4CCE", x"4B756E", x"4B9E02", x"4BC68B", x"4BEF08", x"4C1779", x"4C3FDF", x"4C6839", x"4C9087", x"4CB8C9",
x"4CE0FF", x"4D092A", x"4D3148", x"4D595B", x"4D8162", x"4DA95C", x"4DD14B", x"4DF92E", x"4E2105", x"4E48D0",
x"4E708E", x"4E9841", x"4EBFE8", x"4EE782", x"4F0F10", x"4F3692", x"4F5E08", x"4F8571", x"4FACCF", x"4FD420",
x"4FFB64", x"50229D", x"5049C8", x"5070E8", x"5097FB", x"50BF02", x"50E5FC", x"510CEA", x"5133CB", x"515AA0",
x"518169", x"51A824", x"51CED3", x"51F576", x"521C0C", x"524295", x"526911", x"528F81", x"52B5E4", x"52DC3A",
x"530284", x"5328C1", x"534EF1", x"537514", x"539B2A", x"53C133", x"53E72F", x"540D1F", x"543301", x"5458D7",
x"547E9F", x"54A45B", x"54CA09", x"54EFAA", x"55153F", x"553AC6", x"556040", x"5585AD", x"55AB0C", x"55D05E",
x"55F5A4", x"561ADC", x"564006", x"566523", x"568A33", x"56AF36", x"56D42B", x"56F913", x"571DEE", x"5742BB",
x"57677A", x"578C2D", x"57B0D1", x"57D568", x"57F9F2", x"581E6E", x"5842DC", x"58673D", x"588B90", x"58AFD6",
x"58D40D", x"58F837", x"591C54", x"594063", x"596463", x"598856", x"59AC3C", x"59D013", x"59F3DD", x"5A1799",
x"5A3B46", x"5A5EE6", x"5A8278", x"5AA5FC", x"5AC972", x"5AECDB", x"5B1035", x"5B3381", x"5B56BF", x"5B79EE",
x"5B9D10", x"5BC024", x"5BE329", x"5C0620", x"5C290A", x"5C4BE4", x"5C6EB1", x"5C9170", x"5CB420", x"5CD6C1",
x"5CF955", x"5D1BDA", x"5D3E51", x"5D60B9", x"5D8313", x"5DA55F", x"5DC79C", x"5DE9CB", x"5E0BEB", x"5E2DFD",
x"5E5000", x"5E71F5", x"5E93DB", x"5EB5B2", x"5ED77B", x"5EF936", x"5F1AE1", x"5F3C7E", x"5F5E0C", x"5F7F8C",
x"5FA0FD", x"5FC25F", x"5FE3B2", x"6004F7", x"60262D", x"604753", x"60686C", x"608975", x"60AA6F", x"60CB5A",
x"60EC37", x"610D04", x"612DC3", x"614E73", x"616F13", x"618FA5", x"61B027", x"61D09B", x"61F0FF", x"621154",
x"62319A", x"6251D1", x"6271F9", x"629212", x"62B21B", x"62D215", x"62F200", x"6311DC", x"6331A9", x"635166",
x"637114", x"6390B2", x"63B041", x"63CFC1", x"63EF31", x"640E92", x"642DE4", x"644D26", x"646C58", x"648B7C",
x"64AA8F", x"64C993", x"64E888", x"65076D", x"652642", x"654508", x"6563BE", x"658265", x"65A0FC", x"65BF83",
x"65DDFB", x"65FC62", x"661ABA", x"663903", x"66573B", x"667564", x"66937D", x"66B186", x"66CF80", x"66ED69",
x"670B43", x"67290D", x"6746C7", x"676470", x"67820A", x"679F94", x"67BD0E", x"67DA78", x"67F7D2", x"68151C",
x"683256", x"684F80", x"686C9A", x"6889A4", x"68A69D", x"68C387", x"68E060", x"68FD29", x"6919E2", x"69368A",
x"695323", x"696FAB", x"698C23", x"69A88B", x"69C4E2", x"69E129", x"69FD60", x"6A1986", x"6A359C", x"6A51A2",
x"6A6D97", x"6A897C", x"6AA551", x"6AC115", x"6ADCC8", x"6AF86B", x"6B13FE", x"6B2F80", x"6B4AF1", x"6B6652",
x"6B81A2", x"6B9CE2", x"6BB811", x"6BD330", x"6BEE3E", x"6C093B", x"6C2428", x"6C3F04", x"6C59CF", x"6C748A",
x"6C8F34", x"6CA9CD", x"6CC455", x"6CDECD", x"6CF934", x"6D138A", x"6D2DCF", x"6D4803", x"6D6227", x"6D7C39",
x"6D963B", x"6DB02C", x"6DCA0C", x"6DE3DB", x"6DFD99", x"6E1746", x"6E30E2", x"6E4A6D", x"6E63E7", x"6E7D50",
x"6E96A8", x"6EAFEF", x"6EC925", x"6EE24A", x"6EFB5E", x"6F1460", x"6F2D52", x"6F4632", x"6F5F01", x"6F77BF",
x"6F906C", x"6FA908", x"6FC192", x"6FDA0B", x"6FF273", x"700ACA", x"70230F", x"703B43", x"705366", x"706B78",
x"708378", x"709B66", x"70B344", x"70CB10", x"70E2CA", x"70FA74", x"71120B", x"712992", x"714107", x"71586A",
x"716FBC", x"7186FC", x"719E2B", x"71B549", x"71CC55", x"71E34F", x"71FA38", x"72110F", x"7227D5", x"723E89",
x"72552B", x"726BBC", x"72823B", x"7298A8", x"72AF04", x"72C54E", x"72DB87", x"72F1AD", x"7307C2", x"731DC6",
x"7333B7", x"734997", x"735F65", x"737521", x"738ACB", x"73A064", x"73B5EA", x"73CB5F", x"73E0C2", x"73F613",
x"740B53", x"742080", x"74359B", x"744AA5", x"745F9C", x"747482", x"748956", x"749E17", x"74B2C7", x"74C765",
x"74DBF1", x"74F06A", x"7504D2", x"751927", x"752D6B", x"75419C", x"7555BC", x"7569C9", x"757DC4", x"7591AD",
x"75A584", x"75B949", x"75CCFC", x"75E09C", x"75F42B", x"7607A7", x"761B11", x"762E68", x"7641AE", x"7654E1",
x"766802", x"767B11", x"768E0D", x"76A0F7", x"76B3CF", x"76C695", x"76D948", x"76EBE9", x"76FE78", x"7710F4",
x"77235E", x"7735B5", x"7747FA", x"775A2D", x"776C4D", x"777E5B", x"779057", x"77A240", x"77B416", x"77C5DB",
x"77D78C", x"77E92B", x"77FAB8", x"780C32", x"781D9A", x"782EEF", x"784032", x"785162", x"78627F", x"78738A",
x"788483", x"789568", x"78A63C", x"78B6FC", x"78C7AA", x"78D846", x"78E8CE", x"78F944", x"7909A8", x"7919F8",
x"792A37", x"793A62", x"794A7B", x"795A81", x"796A74", x"797A54", x"798A22", x"7999DD", x"79A986", x"79B91B",
x"79C89E", x"79D80E", x"79E76B", x"79F6B6", x"7A05ED", x"7A1512", x"7A2424", x"7A3323", x"7A420F", x"7A50E9",
x"7A5FAF", x"7A6E63", x"7A7D04", x"7A8B92", x"7A9A0D", x"7AA875", x"7AB6CA", x"7AC50C", x"7AD33C", x"7AE158",
x"7AEF62", x"7AFD58", x"7B0B3C", x"7B190C", x"7B26CA", x"7B3474", x"7B420C", x"7B4F91", x"7B5D02", x"7B6A61",
x"7B77AC", x"7B84E5", x"7B920A", x"7B9F1C", x"7BAC1C", x"7BB908", x"7BC5E1", x"7BD2A7", x"7BDF5A", x"7BEBFA",
x"7BF887", x"7C0500", x"7C1167", x"7C1DBA", x"7C29FA", x"7C3628", x"7C4241", x"7C4E48", x"7C5A3C", x"7C661C",
x"7C71E9", x"7C7DA4", x"7C894A", x"7C94DE", x"7CA05E", x"7CABCC", x"7CB726", x"7CC26C", x"7CCDA0", x"7CD8C0",
x"7CE3CD", x"7CEEC7", x"7CF9AD", x"7D0481", x"7D0F41", x"7D19ED", x"7D2487", x"7D2F0D", x"7D397F", x"7D43DF",
x"7D4E2B", x"7D5864", x"7D6289", x"7D6C9B", x"7D769A", x"7D8086", x"7D8A5E", x"7D9423", x"7D9DD4", x"7DA772",
x"7DB0FC", x"7DBA74", x"7DC3D8", x"7DCD28", x"7DD665", x"7DDF8F", x"7DE8A5", x"7DF1A8", x"7DFA97", x"7E0373",
x"7E0C3C", x"7E14F1", x"7E1D92", x"7E2621", x"7E2E9B", x"7E3703", x"7E3F57", x"7E4797", x"7E4FC4", x"7E57DD",
x"7E5FE3", x"7E67D6", x"7E6FB4", x"7E7780", x"7E7F38", x"7E86DC", x"7E8E6D", x"7E95EB", x"7E9D54", x"7EA4AB",
x"7EABEE", x"7EB31D", x"7EBA39", x"7EC141", x"7EC836", x"7ECF17", x"7ED5E4", x"7EDC9E", x"7EE345", x"7EE9D8",
x"7EF057", x"7EF6C3", x"7EFD1B", x"7F035F", x"7F0990", x"7F0FAE", x"7F15B7", x"7F1BAE", x"7F2190", x"7F275F",
x"7F2D1B", x"7F32C2", x"7F3856", x"7F3DD7", x"7F4344", x"7F489D", x"7F4DE3", x"7F5315", x"7F5833", x"7F5D3E",
x"7F6235", x"7F6719", x"7F6BE8", x"7F70A4", x"7F754D", x"7F79E2", x"7F7E63", x"7F82D1", x"7F872A", x"7F8B71",
x"7F8FA3", x"7F93C2", x"7F97CD", x"7F9BC5", x"7F9FA9", x"7FA379", x"7FA735", x"7FAADE", x"7FAE73", x"7FB1F4",
x"7FB562", x"7FB8BC", x"7FBC03", x"7FBF35", x"7FC254", x"7FC55F", x"7FC857", x"7FCB3B", x"7FCE0B", x"7FD0C7",
x"7FD370", x"7FD605", x"7FD886", x"7FDAF4", x"7FDD4D", x"7FDF94", x"7FE1C6", x"7FE3E5", x"7FE5F0", x"7FE7E7",
x"7FE9CA", x"7FEB9A", x"7FED56", x"7FEEFE", x"7FF093", x"7FF214", x"7FF381", x"7FF4DA", x"7FF620", x"7FF752",
x"7FF870", x"7FF97B", x"7FFA71", x"7FFB54", x"7FFC24", x"7FFCDF", x"7FFD87", x"7FFE1B", x"7FFE9B", x"7FFF08",
x"7FFF61", x"7FFFA6", x"7FFFD7", x"7FFFF5", x"7FFFFF", x"7FFFF5", x"7FFFD7", x"7FFFA6", x"7FFF61", x"7FFF08",
x"7FFE9B", x"7FFE1B", x"7FFD87", x"7FFCDF", x"7FFC24", x"7FFB54", x"7FFA71", x"7FF97B", x"7FF870", x"7FF752",
x"7FF620", x"7FF4DA", x"7FF381", x"7FF214", x"7FF093", x"7FEEFE", x"7FED56", x"7FEB9A", x"7FE9CA", x"7FE7E7",
x"7FE5F0", x"7FE3E5", x"7FE1C6", x"7FDF94", x"7FDD4D", x"7FDAF4", x"7FD886", x"7FD605", x"7FD370", x"7FD0C7",
x"7FCE0B", x"7FCB3B", x"7FC857", x"7FC55F", x"7FC254", x"7FBF35", x"7FBC03", x"7FB8BC", x"7FB562", x"7FB1F4",
x"7FAE73", x"7FAADE", x"7FA735", x"7FA379", x"7F9FA9", x"7F9BC5", x"7F97CD", x"7F93C2", x"7F8FA3", x"7F8B71",
x"7F872A", x"7F82D1", x"7F7E63", x"7F79E2", x"7F754D", x"7F70A4", x"7F6BE8", x"7F6719", x"7F6235", x"7F5D3E",
x"7F5833", x"7F5315", x"7F4DE3", x"7F489D", x"7F4344", x"7F3DD7", x"7F3856", x"7F32C2", x"7F2D1B", x"7F275F",
x"7F2190", x"7F1BAE", x"7F15B7", x"7F0FAE", x"7F0990", x"7F035F", x"7EFD1B", x"7EF6C3", x"7EF057", x"7EE9D8",
x"7EE345", x"7EDC9E", x"7ED5E4", x"7ECF17", x"7EC836", x"7EC141", x"7EBA39", x"7EB31D", x"7EABEE", x"7EA4AB",
x"7E9D54", x"7E95EB", x"7E8E6D", x"7E86DC", x"7E7F38", x"7E7780", x"7E6FB4", x"7E67D6", x"7E5FE3", x"7E57DD",
x"7E4FC4", x"7E4797", x"7E3F57", x"7E3703", x"7E2E9B", x"7E2621", x"7E1D92", x"7E14F1", x"7E0C3C", x"7E0373",
x"7DFA97", x"7DF1A8", x"7DE8A5", x"7DDF8F", x"7DD665", x"7DCD28", x"7DC3D8", x"7DBA74", x"7DB0FC", x"7DA772",
x"7D9DD4", x"7D9423", x"7D8A5E", x"7D8086", x"7D769A", x"7D6C9B", x"7D6289", x"7D5864", x"7D4E2B", x"7D43DF",
x"7D397F", x"7D2F0D", x"7D2487", x"7D19ED", x"7D0F41", x"7D0481", x"7CF9AD", x"7CEEC7", x"7CE3CD", x"7CD8C0",
x"7CCDA0", x"7CC26C", x"7CB726", x"7CABCC", x"7CA05E", x"7C94DE", x"7C894A", x"7C7DA4", x"7C71E9", x"7C661C",
x"7C5A3C", x"7C4E48", x"7C4241", x"7C3628", x"7C29FA", x"7C1DBA", x"7C1167", x"7C0500", x"7BF887", x"7BEBFA",
x"7BDF5A", x"7BD2A7", x"7BC5E1", x"7BB908", x"7BAC1C", x"7B9F1C", x"7B920A", x"7B84E5", x"7B77AC", x"7B6A61",
x"7B5D02", x"7B4F91", x"7B420C", x"7B3474", x"7B26CA", x"7B190C", x"7B0B3C", x"7AFD58", x"7AEF62", x"7AE158",
x"7AD33C", x"7AC50C", x"7AB6CA", x"7AA875", x"7A9A0D", x"7A8B92", x"7A7D04", x"7A6E63", x"7A5FAF", x"7A50E9",
x"7A420F", x"7A3323", x"7A2424", x"7A1512", x"7A05ED", x"79F6B6", x"79E76B", x"79D80E", x"79C89E", x"79B91B",
x"79A986", x"7999DD", x"798A22", x"797A54", x"796A74", x"795A81", x"794A7B", x"793A62", x"792A37", x"7919F8",
x"7909A8", x"78F944", x"78E8CE", x"78D846", x"78C7AA", x"78B6FC", x"78A63C", x"789568", x"788483", x"78738A",
x"78627F", x"785162", x"784032", x"782EEF", x"781D9A", x"780C32", x"77FAB8", x"77E92B", x"77D78C", x"77C5DB",
x"77B416", x"77A240", x"779057", x"777E5B", x"776C4D", x"775A2D", x"7747FA", x"7735B5", x"77235E", x"7710F4",
x"76FE78", x"76EBE9", x"76D948", x"76C695", x"76B3CF", x"76A0F7", x"768E0D", x"767B11", x"766802", x"7654E1",
x"7641AE", x"762E68", x"761B11", x"7607A7", x"75F42B", x"75E09C", x"75CCFC", x"75B949", x"75A584", x"7591AD",
x"757DC4", x"7569C9", x"7555BC", x"75419C", x"752D6B", x"751927", x"7504D2", x"74F06A", x"74DBF1", x"74C765",
x"74B2C7", x"749E17", x"748956", x"747482", x"745F9C", x"744AA5", x"74359B", x"742080", x"740B53", x"73F613",
x"73E0C2", x"73CB5F", x"73B5EA", x"73A064", x"738ACB", x"737521", x"735F65", x"734997", x"7333B7", x"731DC6",
x"7307C2", x"72F1AD", x"72DB87", x"72C54E", x"72AF04", x"7298A8", x"72823B", x"726BBC", x"72552B", x"723E89",
x"7227D5", x"72110F", x"71FA38", x"71E34F", x"71CC55", x"71B549", x"719E2B", x"7186FC", x"716FBC", x"71586A",
x"714107", x"712992", x"71120B", x"70FA74", x"70E2CA", x"70CB10", x"70B344", x"709B66", x"708378", x"706B78",
x"705366", x"703B43", x"70230F", x"700ACA", x"6FF273", x"6FDA0B", x"6FC192", x"6FA908", x"6F906C", x"6F77BF",
x"6F5F01", x"6F4632", x"6F2D52", x"6F1460", x"6EFB5E", x"6EE24A", x"6EC925", x"6EAFEF", x"6E96A8", x"6E7D50",
x"6E63E7", x"6E4A6D", x"6E30E2", x"6E1746", x"6DFD99", x"6DE3DB", x"6DCA0C", x"6DB02C", x"6D963B", x"6D7C39",
x"6D6227", x"6D4803", x"6D2DCF", x"6D138A", x"6CF934", x"6CDECD", x"6CC455", x"6CA9CD", x"6C8F34", x"6C748A",
x"6C59CF", x"6C3F04", x"6C2428", x"6C093B", x"6BEE3E", x"6BD330", x"6BB811", x"6B9CE2", x"6B81A2", x"6B6652",
x"6B4AF1", x"6B2F80", x"6B13FE", x"6AF86B", x"6ADCC8", x"6AC115", x"6AA551", x"6A897C", x"6A6D97", x"6A51A2",
x"6A359C", x"6A1986", x"69FD60", x"69E129", x"69C4E2", x"69A88B", x"698C23", x"696FAB", x"695323", x"69368A",
x"6919E2", x"68FD29", x"68E060", x"68C387", x"68A69D", x"6889A4", x"686C9A", x"684F80", x"683256", x"68151C",
x"67F7D2", x"67DA78", x"67BD0E", x"679F94", x"67820A", x"676470", x"6746C7", x"67290D", x"670B43", x"66ED69",
x"66CF80", x"66B186", x"66937D", x"667564", x"66573B", x"663903", x"661ABA", x"65FC62", x"65DDFB", x"65BF83",
x"65A0FC", x"658265", x"6563BE", x"654508", x"652642", x"65076D", x"64E888", x"64C993", x"64AA8F", x"648B7C",
x"646C58", x"644D26", x"642DE4", x"640E92", x"63EF31", x"63CFC1", x"63B041", x"6390B2", x"637114", x"635166",
x"6331A9", x"6311DC", x"62F200", x"62D215", x"62B21B", x"629212", x"6271F9", x"6251D1", x"62319A", x"621154",
x"61F0FF", x"61D09B", x"61B027", x"618FA5", x"616F13", x"614E73", x"612DC3", x"610D04", x"60EC37", x"60CB5A",
x"60AA6F", x"608975", x"60686C", x"604753", x"60262D", x"6004F7", x"5FE3B2", x"5FC25F", x"5FA0FD", x"5F7F8C",
x"5F5E0C", x"5F3C7E", x"5F1AE1", x"5EF936", x"5ED77B", x"5EB5B2", x"5E93DB", x"5E71F5", x"5E5000", x"5E2DFD",
x"5E0BEB", x"5DE9CB", x"5DC79C", x"5DA55F", x"5D8313", x"5D60B9", x"5D3E51", x"5D1BDA", x"5CF955", x"5CD6C1",
x"5CB420", x"5C9170", x"5C6EB1", x"5C4BE4", x"5C290A", x"5C0620", x"5BE329", x"5BC024", x"5B9D10", x"5B79EE",
x"5B56BF", x"5B3381", x"5B1035", x"5AECDB", x"5AC972", x"5AA5FC", x"5A8278", x"5A5EE6", x"5A3B46", x"5A1799",
x"59F3DD", x"59D013", x"59AC3C", x"598856", x"596463", x"594063", x"591C54", x"58F837", x"58D40D", x"58AFD6",
x"588B90", x"58673D", x"5842DC", x"581E6E", x"57F9F2", x"57D568", x"57B0D1", x"578C2D", x"57677A", x"5742BB",
x"571DEE", x"56F913", x"56D42B", x"56AF36", x"568A33", x"566523", x"564006", x"561ADC", x"55F5A4", x"55D05E",
x"55AB0C", x"5585AD", x"556040", x"553AC6", x"55153F", x"54EFAA", x"54CA09", x"54A45B", x"547E9F", x"5458D7",
x"543301", x"540D1F", x"53E72F", x"53C133", x"539B2A", x"537514", x"534EF1", x"5328C1", x"530284", x"52DC3A",
x"52B5E4", x"528F81", x"526911", x"524295", x"521C0C", x"51F576", x"51CED3", x"51A824", x"518169", x"515AA0",
x"5133CB", x"510CEA", x"50E5FC", x"50BF02", x"5097FB", x"5070E8", x"5049C8", x"50229D", x"4FFB64", x"4FD420",
x"4FACCF", x"4F8571", x"4F5E08", x"4F3692", x"4F0F10", x"4EE782", x"4EBFE8", x"4E9841", x"4E708E", x"4E48D0",
x"4E2105", x"4DF92E", x"4DD14B", x"4DA95C", x"4D8162", x"4D595B", x"4D3148", x"4D092A", x"4CE0FF", x"4CB8C9",
x"4C9087", x"4C6839", x"4C3FDF", x"4C1779", x"4BEF08", x"4BC68B", x"4B9E02", x"4B756E", x"4B4CCE", x"4B2423",
x"4AFB6C", x"4AD2A9", x"4AA9DB", x"4A8101", x"4A581C", x"4A2F2B", x"4A062F", x"49DD27", x"49B414", x"498AF6",
x"4961CC", x"493897", x"490F57", x"48E60B", x"48BCB5", x"489353", x"4869E5", x"48406D", x"4816E9", x"47ED5B",
x"47C3C1", x"479A1C", x"47706D", x"4746B2", x"471CEC", x"46F31B", x"46C93F", x"469F59", x"467567", x"464B6B",
x"462163", x"45F751", x"45CD35", x"45A30D", x"4578DB", x"454E9D", x"452456", x"44FA03", x"44CFA6", x"44A53F",
x"447ACC", x"44504F", x"4425C8", x"43FB36", x"43D09A", x"43A5F3", x"437B42", x"435086", x"4325C0", x"42FAF0",
x"42D015", x"42A530", x"427A41", x"424F47", x"422443", x"41F936", x"41CE1D", x"41A2FB", x"4177CF", x"414C98",
x"412158", x"40F60D", x"40CAB8", x"409F5A", x"4073F1", x"40487F", x"401D02", x"3FF17C", x"3FC5EC", x"3F9A52",
x"3F6EAE", x"3F4300", x"3F1749", x"3EEB88", x"3EBFBD", x"3E93E8", x"3E680A", x"3E3C22", x"3E1031", x"3DE436",
x"3DB832", x"3D8C24", x"3D600C", x"3D33EB", x"3D07C1", x"3CDB8D", x"3CAF50", x"3C8309", x"3C56B9", x"3C2A60",
x"3BFDFE", x"3BD192", x"3BA51D", x"3B789F", x"3B4C18", x"3B1F87", x"3AF2EE", x"3AC64B", x"3A999F", x"3A6CEB",
x"3A402D", x"3A1366", x"39E696", x"39B9BE", x"398CDC", x"395FF2", x"3932FF", x"390603", x"38D8FE", x"38ABF0",
x"387EDA", x"3851BB", x"382493", x"37F762", x"37CA29", x"379CE8", x"376F9D", x"37424B", x"3714EF", x"36E78B",
x"36BA1F", x"368CAA", x"365F2D", x"3631A8", x"36041A", x"35D684", x"35A8E5", x"357B3E", x"354D8F", x"351FD8",
x"34F219", x"34C451", x"349681", x"3468AA", x"343ACA", x"340CE2", x"33DEF2", x"33B0FA", x"3382FA", x"3354F2",
x"3326E2", x"32F8CA", x"32CAAB", x"329C83", x"326E54", x"32401D", x"3211DE", x"31E398", x"31B549", x"3186F4",
x"315896", x"312A31", x"30FBC4", x"30CD50", x"309ED4", x"307051", x"3041C7", x"301334", x"2FE49B", x"2FB5FA",
x"2F8752", x"2F58A2", x"2F29EB", x"2EFB2D", x"2ECC67", x"2E9D9B", x"2E6EC7", x"2E3FEC", x"2E110A", x"2DE220",
x"2DB330", x"2D8439", x"2D553A", x"2D2635", x"2CF728", x"2CC815", x"2C98FB", x"2C69DA", x"2C3AB2", x"2C0B83",
x"2BDC4E", x"2BAD11", x"2B7DCE", x"2B4E85", x"2B1F34", x"2AEFDD", x"2AC07F", x"2A911B", x"2A61B0", x"2A323F",
x"2A02C7", x"29D349", x"29A3C4", x"297438", x"2944A7", x"29150F", x"28E570", x"28B5CC", x"288621", x"285670",
x"2826B8", x"27F6FB", x"27C737", x"27976D", x"27679D", x"2737C7", x"2707EB", x"26D809", x"26A821", x"267833",
x"26483F", x"261845", x"25E845", x"25B83F", x"258834", x"255823", x"25280C", x"24F7EF", x"24C7CC", x"2497A4",
x"246777", x"243743", x"24070A", x"23D6CC", x"23A688", x"23763E", x"2345EF", x"23159B", x"22E541", x"22B4E2",
x"22847D", x"225413", x"2223A4", x"21F330", x"21C2B6", x"219237", x"2161B3", x"21312A", x"21009B", x"20D008",
x"209F6F", x"206ED2", x"203E2F", x"200D88", x"1FDCDB", x"1FAC2A", x"1F7B74", x"1F4AB9", x"1F19F9", x"1EE934",
x"1EB86B", x"1E879C", x"1E56C9", x"1E25F2", x"1DF516", x"1DC435", x"1D934F", x"1D6265", x"1D3177", x"1D0084",
x"1CCF8C", x"1C9E90", x"1C6D90", x"1C3C8B", x"1C0B82", x"1BDA74", x"1BA962", x"1B784C", x"1B4732", x"1B1614",
x"1AE4F1", x"1AB3CA", x"1A829F", x"1A5170", x"1A203D", x"19EF06", x"19BDCB", x"198C8C", x"195B49", x"192A02",
x"18F8B8", x"18C769", x"189616", x"1864C0", x"183366", x"180208", x"17D0A7", x"179F42", x"176DD9", x"173C6D",
x"170AFD", x"16D989", x"16A812", x"167698", x"16451A", x"161398", x"15E214", x"15B08B", x"157F00", x"154D71",
x"151BDF", x"14EA49", x"14B8B1", x"148715", x"145576", x"1423D4", x"13F22F", x"13C086", x"138EDB", x"135D2D",
x"132B7B", x"12F9C7", x"12C810", x"129656", x"126499", x"1232D9", x"120116", x"11CF51", x"119D89", x"116BBE",
x"1139F0", x"110820", x"10D64D", x"10A478", x"1072A0", x"1040C5", x"100EE8", x"0FDD09", x"0FAB27", x"0F7942",
x"0F475B", x"0F1572", x"0EE387", x"0EB199", x"0E7FA9", x"0E4DB7", x"0E1BC2", x"0DE9CC", x"0DB7D3", x"0D85D8",
x"0D53DB", x"0D21DC", x"0CEFDB", x"0CBDD8", x"0C8BD3", x"0C59CC", x"0C27C3", x"0BF5B8", x"0BC3AC", x"0B919D",
x"0B5F8D", x"0B2D7B", x"0AFB67", x"0AC952", x"0A973B", x"0A6522", x"0A3308", x"0A00EC", x"09CECF", x"099CB0",
x"096A90", x"09386E", x"09064B", x"08D426", x"08A200", x"086FD9", x"083DB0", x"080B86", x"07D95B", x"07A72F",
x"077501", x"0742D3", x"0710A3", x"06DE72", x"06AC40", x"067A0D", x"0647D9", x"0615A4", x"05E36E", x"05B137",
x"057F00", x"054CC7", x"051A8E", x"04E854", x"04B619", x"0483DD", x"0451A1", x"041F64", x"03ED26", x"03BAE8",
x"0388A9", x"03566A", x"03242A", x"02F1EA", x"02BFA9", x"028D68", x"025B26", x"0228E4", x"01F6A2", x"01C45F",
x"01921D", x"015FDA", x"012D96", x"00FB53", x"00C90F", x"0096CB", x"006487", x"003243", x"000000", x"FFCDBD",
x"FF9B79", x"FF6935", x"FF36F1", x"FF04AD", x"FED26A", x"FEA026", x"FE6DE3", x"FE3BA1", x"FE095E", x"FDD71C",
x"FDA4DA", x"FD7298", x"FD4057", x"FD0E16", x"FCDBD6", x"FCA996", x"FC7757", x"FC4518", x"FC12DA", x"FBE09C",
x"FBAE5F", x"FB7C23", x"FB49E7", x"FB17AC", x"FAE572", x"FAB339", x"FA8100", x"FA4EC9", x"FA1C92", x"F9EA5C",
x"F9B827", x"F985F3", x"F953C0", x"F9218E", x"F8EF5D", x"F8BD2D", x"F88AFF", x"F858D1", x"F826A5", x"F7F47A",
x"F7C250", x"F79027", x"F75E00", x"F72BDA", x"F6F9B5", x"F6C792", x"F69570", x"F66350", x"F63131", x"F5FF14",
x"F5CCF8", x"F59ADE", x"F568C5", x"F536AE", x"F50499", x"F4D285", x"F4A073", x"F46E63", x"F43C54", x"F40A48",
x"F3D83D", x"F3A634", x"F3742D", x"F34228", x"F31025", x"F2DE24", x"F2AC25", x"F27A28", x"F2482D", x"F21634",
x"F1E43E", x"F1B249", x"F18057", x"F14E67", x"F11C79", x"F0EA8E", x"F0B8A5", x"F086BE", x"F054D9", x"F022F7",
x"EFF118", x"EFBF3B", x"EF8D60", x"EF5B88", x"EF29B3", x"EEF7E0", x"EEC610", x"EE9442", x"EE6277", x"EE30AF",
x"EDFEEA", x"EDCD27", x"ED9B67", x"ED69AA", x"ED37F0", x"ED0639", x"ECD485", x"ECA2D3", x"EC7125", x"EC3F7A",
x"EC0DD1", x"EBDC2C", x"EBAA8A", x"EB78EB", x"EB474F", x"EB15B7", x"EAE421", x"EAB28F", x"EA8100", x"EA4F75",
x"EA1DEC", x"E9EC68", x"E9BAE6", x"E98968", x"E957EE", x"E92677", x"E8F503", x"E8C393", x"E89227", x"E860BE",
x"E82F59", x"E7FDF8", x"E7CC9A", x"E79B40", x"E769EA", x"E73897", x"E70748", x"E6D5FE", x"E6A4B7", x"E67374",
x"E64235", x"E610FA", x"E5DFC3", x"E5AE90", x"E57D61", x"E54C36", x"E51B0F", x"E4E9EC", x"E4B8CE", x"E487B4",
x"E4569E", x"E4258C", x"E3F47E", x"E3C375", x"E39270", x"E36170", x"E33074", x"E2FF7C", x"E2CE89", x"E29D9B",
x"E26CB1", x"E23BCB", x"E20AEA", x"E1DA0E", x"E1A937", x"E17864", x"E14795", x"E116CC", x"E0E607", x"E0B547",
x"E0848C", x"E053D6", x"E02325", x"DFF278", x"DFC1D1", x"DF912E", x"DF6091", x"DF2FF8", x"DEFF65", x"DECED6",
x"DE9E4D", x"DE6DC9", x"DE3D4A", x"DE0CD0", x"DDDC5C", x"DDABED", x"DD7B83", x"DD4B1E", x"DD1ABF", x"DCEA65",
x"DCBA11", x"DC89C2", x"DC5978", x"DC2934", x"DBF8F6", x"DBC8BD", x"DB9889", x"DB685C", x"DB3834", x"DB0811",
x"DAD7F4", x"DAA7DD", x"DA77CC", x"DA47C1", x"DA17BB", x"D9E7BB", x"D9B7C1", x"D987CD", x"D957DF", x"D927F7",
x"D8F815", x"D8C839", x"D89863", x"D86893", x"D838C9", x"D80905", x"D7D948", x"D7A990", x"D779DF", x"D74A34",
x"D71A90", x"D6EAF1", x"D6BB59", x"D68BC8", x"D65C3C", x"D62CB7", x"D5FD39", x"D5CDC1", x"D59E50", x"D56EE5",
x"D53F81", x"D51023", x"D4E0CC", x"D4B17B", x"D48232", x"D452EF", x"D423B2", x"D3F47D", x"D3C54E", x"D39626",
x"D36705", x"D337EB", x"D308D8", x"D2D9CB", x"D2AAC6", x"D27BC7", x"D24CD0", x"D21DE0", x"D1EEF6", x"D1C014",
x"D19139", x"D16265", x"D13399", x"D104D3", x"D0D615", x"D0A75E", x"D078AE", x"D04A06", x"D01B65", x"CFECCC",
x"CFBE39", x"CF8FAF", x"CF612C", x"CF32B0", x"CF043C", x"CED5CF", x"CEA76A", x"CE790C", x"CE4AB7", x"CE1C68",
x"CDEE22", x"CDBFE3", x"CD91AC", x"CD637D", x"CD3555", x"CD0736", x"CCD91E", x"CCAB0E", x"CC7D06", x"CC4F06",
x"CC210E", x"CBF31E", x"CBC536", x"CB9756", x"CB697F", x"CB3BAF", x"CB0DE7", x"CAE028", x"CAB271", x"CA84C2",
x"CA571B", x"CA297C", x"C9FBE6", x"C9CE58", x"C9A0D3", x"C97356", x"C945E1", x"C91875", x"C8EB11", x"C8BDB5",
x"C89063", x"C86318", x"C835D7", x"C8089E", x"C7DB6D", x"C7AE45", x"C78126", x"C75410", x"C72702", x"C6F9FD",
x"C6CD01", x"C6A00E", x"C67324", x"C64642", x"C6196A", x"C5EC9A", x"C5BFD3", x"C59315", x"C56661", x"C539B5",
x"C50D12", x"C4E079", x"C4B3E8", x"C48761", x"C45AE3", x"C42E6E", x"C40202", x"C3D5A0", x"C3A947", x"C37CF7",
x"C350B0", x"C32473", x"C2F83F", x"C2CC15", x"C29FF4", x"C273DC", x"C247CE", x"C21BCA", x"C1EFCF", x"C1C3DE",
x"C197F6", x"C16C18", x"C14043", x"C11478", x"C0E8B7", x"C0BD00", x"C09152", x"C065AE", x"C03A14", x"C00E84",
x"BFE2FE", x"BFB781", x"BF8C0F", x"BF60A6", x"BF3548", x"BF09F3", x"BEDEA8", x"BEB368", x"BE8831", x"BE5D05",
x"BE31E3", x"BE06CA", x"BDDBBD", x"BDB0B9", x"BD85BF", x"BD5AD0", x"BD2FEB", x"BD0510", x"BCDA40", x"BCAF7A",
x"BC84BE", x"BC5A0D", x"BC2F66", x"BC04CA", x"BBDA38", x"BBAFB1", x"BB8534", x"BB5AC1", x"BB305A", x"BB05FD",
x"BADBAA", x"BAB163", x"BA8725", x"BA5CF3", x"BA32CB", x"BA08AF", x"B9DE9D", x"B9B495", x"B98A99", x"B960A7",
x"B936C1", x"B90CE5", x"B8E314", x"B8B94E", x"B88F93", x"B865E4", x"B83C3F", x"B812A5", x"B7E917", x"B7BF93",
x"B7961B", x"B76CAD", x"B7434B", x"B719F5", x"B6F0A9", x"B6C769", x"B69E34", x"B6750A", x"B64BEC", x"B622D9",
x"B5F9D1", x"B5D0D5", x"B5A7E4", x"B57EFF", x"B55625", x"B52D57", x"B50494", x"B4DBDD", x"B4B332", x"B48A92",
x"B461FE", x"B43975", x"B410F8", x"B3E887", x"B3C021", x"B397C7", x"B36F79", x"B34737", x"B31F01", x"B2F6D6",
x"B2CEB8", x"B2A6A5", x"B27E9E", x"B256A4", x"B22EB5", x"B206D2", x"B1DEFB", x"B1B730", x"B18F72", x"B167BF",
x"B14018", x"B1187E", x"B0F0F0", x"B0C96E", x"B0A1F8", x"B07A8F", x"B05331", x"B02BE0", x"B0049C", x"AFDD63",
x"AFB638", x"AF8F18", x"AF6805", x"AF40FE", x"AF1A04", x"AEF316", x"AECC35", x"AEA560", x"AE7E97", x"AE57DC",
x"AE312D", x"AE0A8A", x"ADE3F4", x"ADBD6B", x"AD96EF", x"AD707F", x"AD4A1C", x"AD23C6", x"ACFD7C", x"ACD73F",
x"ACB10F", x"AC8AEC", x"AC64D6", x"AC3ECD", x"AC18D1", x"ABF2E1", x"ABCCFF", x"ABA729", x"AB8161", x"AB5BA5",
x"AB35F7", x"AB1056", x"AAEAC1", x"AAC53A", x"AA9FC0", x"AA7A53", x"AA54F4", x"AA2FA2", x"AA0A5C", x"A9E524",
x"A9BFFA", x"A99ADD", x"A975CD", x"A950CA", x"A92BD5", x"A906ED", x"A8E212", x"A8BD45", x"A89886", x"A873D3",
x"A84F2F", x"A82A98", x"A8060E", x"A7E192", x"A7BD24", x"A798C3", x"A77470", x"A7502A", x"A72BF3", x"A707C9",
x"A6E3AC", x"A6BF9D", x"A69B9D", x"A677AA", x"A653C4", x"A62FED", x"A60C23", x"A5E867", x"A5C4BA", x"A5A11A",
x"A57D88", x"A55A04", x"A5368E", x"A51325", x"A4EFCB", x"A4CC7F", x"A4A941", x"A48612", x"A462F0", x"A43FDC",
x"A41CD7", x"A3F9E0", x"A3D6F6", x"A3B41C", x"A3914F", x"A36E90", x"A34BE0", x"A3293F", x"A306AB", x"A2E426",
x"A2C1AF", x"A29F47", x"A27CED", x"A25AA1", x"A23864", x"A21635", x"A1F415", x"A1D203", x"A1B000", x"A18E0B",
x"A16C25", x"A14A4E", x"A12885", x"A106CA", x"A0E51F", x"A0C382", x"A0A1F4", x"A08074", x"A05F03", x"A03DA1",
x"A01C4E", x"9FFB09", x"9FD9D3", x"9FB8AD", x"9F9794", x"9F768B", x"9F5591", x"9F34A6", x"9F13C9", x"9EF2FC",
x"9ED23D", x"9EB18D", x"9E90ED", x"9E705B", x"9E4FD9", x"9E2F65", x"9E0F01", x"9DEEAC", x"9DCE66", x"9DAE2F",
x"9D8E07", x"9D6DEE", x"9D4DE5", x"9D2DEB", x"9D0E00", x"9CEE24", x"9CCE57", x"9CAE9A", x"9C8EEC", x"9C6F4E",
x"9C4FBF", x"9C303F", x"9C10CF", x"9BF16E", x"9BD21C", x"9BB2DA", x"9B93A8", x"9B7484", x"9B5571", x"9B366D",
x"9B1778", x"9AF893", x"9AD9BE", x"9ABAF8", x"9A9C42", x"9A7D9B", x"9A5F04", x"9A407D", x"9A2205", x"9A039E",
x"99E546", x"99C6FD", x"99A8C5", x"998A9C", x"996C83", x"994E7A", x"993080", x"991297", x"98F4BD", x"98D6F3",
x"98B939", x"989B90", x"987DF6", x"98606C", x"9842F2", x"982588", x"98082E", x"97EAE4", x"97CDAA", x"97B080",
x"979366", x"97765C", x"975963", x"973C79", x"971FA0", x"9702D7", x"96E61E", x"96C976", x"96ACDD", x"969055",
x"9673DD", x"965775", x"963B1E", x"961ED7", x"9602A0", x"95E67A", x"95CA64", x"95AE5E", x"959269", x"957684",
x"955AAF", x"953EEB", x"952338", x"950795", x"94EC02", x"94D080", x"94B50F", x"9499AE", x"947E5E", x"94631E",
x"9447EF", x"942CD0", x"9411C2", x"93F6C5", x"93DBD8", x"93C0FC", x"93A631", x"938B76", x"9370CC", x"935633",
x"933BAB", x"932133", x"9306CC", x"92EC76", x"92D231", x"92B7FD", x"929DD9", x"9283C7", x"9269C5", x"924FD4",
x"9235F4", x"921C25", x"920267", x"91E8BA", x"91CF1E", x"91B593", x"919C19", x"9182B0", x"916958", x"915011",
x"9136DB", x"911DB6", x"9104A2", x"90EBA0", x"90D2AE", x"90B9CE", x"90A0FF", x"908841", x"906F94", x"9056F8",
x"903E6E", x"9025F5", x"900D8D", x"8FF536", x"8FDCF1", x"8FC4BD", x"8FAC9A", x"8F9488", x"8F7C88", x"8F649A",
x"8F4CBC", x"8F34F0", x"8F1D36", x"8F058C", x"8EEDF5", x"8ED66E", x"8EBEF9", x"8EA796", x"8E9044", x"8E7904",
x"8E61D5", x"8E4AB7", x"8E33AB", x"8E1CB1", x"8E05C8", x"8DEEF1", x"8DD82B", x"8DC177", x"8DAAD5", x"8D9444",
x"8D7DC5", x"8D6758", x"8D50FC", x"8D3AB2", x"8D2479", x"8D0E53", x"8CF83E", x"8CE23A", x"8CCC49", x"8CB669",
x"8CA09B", x"8C8ADF", x"8C7535", x"8C5F9C", x"8C4A16", x"8C34A1", x"8C1F3E", x"8C09ED", x"8BF4AD", x"8BDF80",
x"8BCA65", x"8BB55B", x"8BA064", x"8B8B7E", x"8B76AA", x"8B61E9", x"8B4D39", x"8B389B", x"8B240F", x"8B0F96",
x"8AFB2E", x"8AE6D9", x"8AD295", x"8ABE64", x"8AAA44", x"8A9637", x"8A823C", x"8A6E53", x"8A5A7C", x"8A46B7",
x"8A3304", x"8A1F64", x"8A0BD5", x"89F859", x"89E4EF", x"89D198", x"89BE52", x"89AB1F", x"8997FE", x"8984EF",
x"8971F3", x"895F09", x"894C31", x"89396B", x"8926B8", x"891417", x"890188", x"88EF0C", x"88DCA2", x"88CA4B",
x"88B806", x"88A5D3", x"8893B3", x"8881A5", x"886FA9", x"885DC0", x"884BEA", x"883A25", x"882874", x"8816D5",
x"880548", x"87F3CE", x"87E266", x"87D111", x"87BFCE", x"87AE9E", x"879D81", x"878C76", x"877B7D", x"876A98",
x"8759C4", x"874904", x"873856", x"8727BA", x"871732", x"8706BC", x"86F658", x"86E608", x"86D5C9", x"86C59E",
x"86B585", x"86A57F", x"86958C", x"8685AC", x"8675DE", x"866623", x"86567A", x"8646E5", x"863762", x"8627F2",
x"861895", x"86094A", x"85FA13", x"85EAEE", x"85DBDC", x"85CCDD", x"85BDF1", x"85AF17", x"85A051", x"85919D",
x"8582FC", x"85746E", x"8565F3", x"85578B", x"854936", x"853AF4", x"852CC4", x"851EA8", x"85109E", x"8502A8",
x"84F4C4", x"84E6F4", x"84D936", x"84CB8C", x"84BDF4", x"84B06F", x"84A2FE", x"84959F", x"848854", x"847B1B",
x"846DF6", x"8460E4", x"8453E4", x"8446F8", x"843A1F", x"842D59", x"8420A6", x"841406", x"840779", x"83FB00",
x"83EE99", x"83E246", x"83D606", x"83C9D8", x"83BDBF", x"83B1B8", x"83A5C4", x"8399E4", x"838E17", x"83825C",
x"8376B6", x"836B22", x"835FA2", x"835434", x"8348DA", x"833D94", x"833260", x"832740", x"831C33", x"831139",
x"830653", x"82FB7F", x"82F0BF", x"82E613", x"82DB79", x"82D0F3", x"82C681", x"82BC21", x"82B1D5", x"82A79C",
x"829D77", x"829365", x"828966", x"827F7A", x"8275A2", x"826BDD", x"82622C", x"82588E", x"824F04", x"82458C",
x"823C28", x"8232D8", x"82299B", x"822071", x"82175B", x"820E58", x"820569", x"81FC8D", x"81F3C4", x"81EB0F",
x"81E26E", x"81D9DF", x"81D165", x"81C8FD", x"81C0A9", x"81B869", x"81B03C", x"81A823", x"81A01D", x"81982A",
x"81904C", x"818880", x"8180C8", x"817924", x"817193", x"816A15", x"8162AC", x"815B55", x"815412", x"814CE3",
x"8145C7", x"813EBF", x"8137CA", x"8130E9", x"812A1C", x"812362", x"811CBB", x"811628", x"810FA9", x"81093D",
x"8102E5", x"80FCA1", x"80F670", x"80F052", x"80EA49", x"80E452", x"80DE70", x"80D8A1", x"80D2E5", x"80CD3E",
x"80C7AA", x"80C229", x"80BCBC", x"80B763", x"80B21D", x"80ACEB", x"80A7CD", x"80A2C2", x"809DCB", x"8098E7",
x"809418", x"808F5C", x"808AB3", x"80861E", x"80819D", x"807D2F", x"8078D6", x"80748F", x"80705D", x"806C3E",
x"806833", x"80643B", x"806057", x"805C87", x"8058CB", x"805522", x"80518D", x"804E0C", x"804A9E", x"804744",
x"8043FD", x"8040CB", x"803DAC", x"803AA1", x"8037A9", x"8034C5", x"8031F5", x"802F39", x"802C90", x"8029FB",
x"80277A", x"80250C", x"8022B3", x"80206C", x"801E3A", x"801C1B", x"801A10", x"801819", x"801636", x"801466",
x"8012AA", x"801102", x"800F6D", x"800DEC", x"800C7F", x"800B26", x"8009E0", x"8008AE", x"800790", x"800685",
x"80058F", x"8004AC", x"8003DC", x"800321", x"800279", x"8001E5", x"800165", x"8000F8", x"80009F", x"80005A",
x"800029", x"80000B", x"800001", x"80000B", x"800029", x"80005A", x"80009F", x"8000F8", x"800165", x"8001E5",
x"800279", x"800321", x"8003DC", x"8004AC", x"80058F", x"800685", x"800790", x"8008AE", x"8009E0", x"800B26",
x"800C7F", x"800DEC", x"800F6D", x"801102", x"8012AA", x"801466", x"801636", x"801819", x"801A10", x"801C1B",
x"801E3A", x"80206C", x"8022B3", x"80250C", x"80277A", x"8029FB", x"802C90", x"802F39", x"8031F5", x"8034C5",
x"8037A9", x"803AA1", x"803DAC", x"8040CB", x"8043FD", x"804744", x"804A9E", x"804E0C", x"80518D", x"805522",
x"8058CB", x"805C87", x"806057", x"80643B", x"806833", x"806C3E", x"80705D", x"80748F", x"8078D6", x"807D2F",
x"80819D", x"80861E", x"808AB3", x"808F5C", x"809418", x"8098E7", x"809DCB", x"80A2C2", x"80A7CD", x"80ACEB",
x"80B21D", x"80B763", x"80BCBC", x"80C229", x"80C7AA", x"80CD3E", x"80D2E5", x"80D8A1", x"80DE70", x"80E452",
x"80EA49", x"80F052", x"80F670", x"80FCA1", x"8102E5", x"81093D", x"810FA9", x"811628", x"811CBB", x"812362",
x"812A1C", x"8130E9", x"8137CA", x"813EBF", x"8145C7", x"814CE3", x"815412", x"815B55", x"8162AC", x"816A15",
x"817193", x"817924", x"8180C8", x"818880", x"81904C", x"81982A", x"81A01D", x"81A823", x"81B03C", x"81B869",
x"81C0A9", x"81C8FD", x"81D165", x"81D9DF", x"81E26E", x"81EB0F", x"81F3C4", x"81FC8D", x"820569", x"820E58",
x"82175B", x"822071", x"82299B", x"8232D8", x"823C28", x"82458C", x"824F04", x"82588E", x"82622C", x"826BDD",
x"8275A2", x"827F7A", x"828966", x"829365", x"829D77", x"82A79C", x"82B1D5", x"82BC21", x"82C681", x"82D0F3",
x"82DB79", x"82E613", x"82F0BF", x"82FB7F", x"830653", x"831139", x"831C33", x"832740", x"833260", x"833D94",
x"8348DA", x"835434", x"835FA2", x"836B22", x"8376B6", x"83825C", x"838E17", x"8399E4", x"83A5C4", x"83B1B8",
x"83BDBF", x"83C9D8", x"83D606", x"83E246", x"83EE99", x"83FB00", x"840779", x"841406", x"8420A6", x"842D59",
x"843A1F", x"8446F8", x"8453E4", x"8460E4", x"846DF6", x"847B1B", x"848854", x"84959F", x"84A2FE", x"84B06F",
x"84BDF4", x"84CB8C", x"84D936", x"84E6F4", x"84F4C4", x"8502A8", x"85109E", x"851EA8", x"852CC4", x"853AF4",
x"854936", x"85578B", x"8565F3", x"85746E", x"8582FC", x"85919D", x"85A051", x"85AF17", x"85BDF1", x"85CCDD",
x"85DBDC", x"85EAEE", x"85FA13", x"86094A", x"861895", x"8627F2", x"863762", x"8646E5", x"86567A", x"866623",
x"8675DE", x"8685AC", x"86958C", x"86A57F", x"86B585", x"86C59E", x"86D5C9", x"86E608", x"86F658", x"8706BC",
x"871732", x"8727BA", x"873856", x"874904", x"8759C4", x"876A98", x"877B7D", x"878C76", x"879D81", x"87AE9E",
x"87BFCE", x"87D111", x"87E266", x"87F3CE", x"880548", x"8816D5", x"882874", x"883A25", x"884BEA", x"885DC0",
x"886FA9", x"8881A5", x"8893B3", x"88A5D3", x"88B806", x"88CA4B", x"88DCA2", x"88EF0C", x"890188", x"891417",
x"8926B8", x"89396B", x"894C31", x"895F09", x"8971F3", x"8984EF", x"8997FE", x"89AB1F", x"89BE52", x"89D198",
x"89E4EF", x"89F859", x"8A0BD5", x"8A1F64", x"8A3304", x"8A46B7", x"8A5A7C", x"8A6E53", x"8A823C", x"8A9637",
x"8AAA44", x"8ABE64", x"8AD295", x"8AE6D9", x"8AFB2E", x"8B0F96", x"8B240F", x"8B389B", x"8B4D39", x"8B61E9",
x"8B76AA", x"8B8B7E", x"8BA064", x"8BB55B", x"8BCA65", x"8BDF80", x"8BF4AD", x"8C09ED", x"8C1F3E", x"8C34A1",
x"8C4A16", x"8C5F9C", x"8C7535", x"8C8ADF", x"8CA09B", x"8CB669", x"8CCC49", x"8CE23A", x"8CF83E", x"8D0E53",
x"8D2479", x"8D3AB2", x"8D50FC", x"8D6758", x"8D7DC5", x"8D9444", x"8DAAD5", x"8DC177", x"8DD82B", x"8DEEF1",
x"8E05C8", x"8E1CB1", x"8E33AB", x"8E4AB7", x"8E61D5", x"8E7904", x"8E9044", x"8EA796", x"8EBEF9", x"8ED66E",
x"8EEDF5", x"8F058C", x"8F1D36", x"8F34F0", x"8F4CBC", x"8F649A", x"8F7C88", x"8F9488", x"8FAC9A", x"8FC4BD",
x"8FDCF1", x"8FF536", x"900D8D", x"9025F5", x"903E6E", x"9056F8", x"906F94", x"908841", x"90A0FF", x"90B9CE",
x"90D2AE", x"90EBA0", x"9104A2", x"911DB6", x"9136DB", x"915011", x"916958", x"9182B0", x"919C19", x"91B593",
x"91CF1E", x"91E8BA", x"920267", x"921C25", x"9235F4", x"924FD4", x"9269C5", x"9283C7", x"929DD9", x"92B7FD",
x"92D231", x"92EC76", x"9306CC", x"932133", x"933BAB", x"935633", x"9370CC", x"938B76", x"93A631", x"93C0FC",
x"93DBD8", x"93F6C5", x"9411C2", x"942CD0", x"9447EF", x"94631E", x"947E5E", x"9499AE", x"94B50F", x"94D080",
x"94EC02", x"950795", x"952338", x"953EEB", x"955AAF", x"957684", x"959269", x"95AE5E", x"95CA64", x"95E67A",
x"9602A0", x"961ED7", x"963B1E", x"965775", x"9673DD", x"969055", x"96ACDD", x"96C976", x"96E61E", x"9702D7",
x"971FA0", x"973C79", x"975963", x"97765C", x"979366", x"97B080", x"97CDAA", x"97EAE4", x"98082E", x"982588",
x"9842F2", x"98606C", x"987DF6", x"989B90", x"98B939", x"98D6F3", x"98F4BD", x"991297", x"993080", x"994E7A",
x"996C83", x"998A9C", x"99A8C5", x"99C6FD", x"99E546", x"9A039E", x"9A2205", x"9A407D", x"9A5F04", x"9A7D9B",
x"9A9C42", x"9ABAF8", x"9AD9BE", x"9AF893", x"9B1778", x"9B366D", x"9B5571", x"9B7484", x"9B93A8", x"9BB2DA",
x"9BD21C", x"9BF16E", x"9C10CF", x"9C303F", x"9C4FBF", x"9C6F4E", x"9C8EEC", x"9CAE9A", x"9CCE57", x"9CEE24",
x"9D0E00", x"9D2DEB", x"9D4DE5", x"9D6DEE", x"9D8E07", x"9DAE2F", x"9DCE66", x"9DEEAC", x"9E0F01", x"9E2F65",
x"9E4FD9", x"9E705B", x"9E90ED", x"9EB18D", x"9ED23D", x"9EF2FC", x"9F13C9", x"9F34A6", x"9F5591", x"9F768B",
x"9F9794", x"9FB8AD", x"9FD9D3", x"9FFB09", x"A01C4E", x"A03DA1", x"A05F03", x"A08074", x"A0A1F4", x"A0C382",
x"A0E51F", x"A106CA", x"A12885", x"A14A4E", x"A16C25", x"A18E0B", x"A1B000", x"A1D203", x"A1F415", x"A21635",
x"A23864", x"A25AA1", x"A27CED", x"A29F47", x"A2C1AF", x"A2E426", x"A306AB", x"A3293F", x"A34BE0", x"A36E90",
x"A3914F", x"A3B41C", x"A3D6F6", x"A3F9E0", x"A41CD7", x"A43FDC", x"A462F0", x"A48612", x"A4A941", x"A4CC7F",
x"A4EFCB", x"A51325", x"A5368E", x"A55A04", x"A57D88", x"A5A11A", x"A5C4BA", x"A5E867", x"A60C23", x"A62FED",
x"A653C4", x"A677AA", x"A69B9D", x"A6BF9D", x"A6E3AC", x"A707C9", x"A72BF3", x"A7502A", x"A77470", x"A798C3",
x"A7BD24", x"A7E192", x"A8060E", x"A82A98", x"A84F2F", x"A873D3", x"A89886", x"A8BD45", x"A8E212", x"A906ED",
x"A92BD5", x"A950CA", x"A975CD", x"A99ADD", x"A9BFFA", x"A9E524", x"AA0A5C", x"AA2FA2", x"AA54F4", x"AA7A53",
x"AA9FC0", x"AAC53A", x"AAEAC1", x"AB1056", x"AB35F7", x"AB5BA5", x"AB8161", x"ABA729", x"ABCCFF", x"ABF2E1",
x"AC18D1", x"AC3ECD", x"AC64D6", x"AC8AEC", x"ACB10F", x"ACD73F", x"ACFD7C", x"AD23C6", x"AD4A1C", x"AD707F",
x"AD96EF", x"ADBD6B", x"ADE3F4", x"AE0A8A", x"AE312D", x"AE57DC", x"AE7E97", x"AEA560", x"AECC35", x"AEF316",
x"AF1A04", x"AF40FE", x"AF6805", x"AF8F18", x"AFB638", x"AFDD63", x"B0049C", x"B02BE0", x"B05331", x"B07A8F",
x"B0A1F8", x"B0C96E", x"B0F0F0", x"B1187E", x"B14018", x"B167BF", x"B18F72", x"B1B730", x"B1DEFB", x"B206D2",
x"B22EB5", x"B256A4", x"B27E9E", x"B2A6A5", x"B2CEB8", x"B2F6D6", x"B31F01", x"B34737", x"B36F79", x"B397C7",
x"B3C021", x"B3E887", x"B410F8", x"B43975", x"B461FE", x"B48A92", x"B4B332", x"B4DBDD", x"B50494", x"B52D57",
x"B55625", x"B57EFF", x"B5A7E4", x"B5D0D5", x"B5F9D1", x"B622D9", x"B64BEC", x"B6750A", x"B69E34", x"B6C769",
x"B6F0A9", x"B719F5", x"B7434B", x"B76CAD", x"B7961B", x"B7BF93", x"B7E917", x"B812A5", x"B83C3F", x"B865E4",
x"B88F93", x"B8B94E", x"B8E314", x"B90CE5", x"B936C1", x"B960A7", x"B98A99", x"B9B495", x"B9DE9D", x"BA08AF",
x"BA32CB", x"BA5CF3", x"BA8725", x"BAB163", x"BADBAA", x"BB05FD", x"BB305A", x"BB5AC1", x"BB8534", x"BBAFB1",
x"BBDA38", x"BC04CA", x"BC2F66", x"BC5A0D", x"BC84BE", x"BCAF7A", x"BCDA40", x"BD0510", x"BD2FEB", x"BD5AD0",
x"BD85BF", x"BDB0B9", x"BDDBBD", x"BE06CA", x"BE31E3", x"BE5D05", x"BE8831", x"BEB368", x"BEDEA8", x"BF09F3",
x"BF3548", x"BF60A6", x"BF8C0F", x"BFB781", x"BFE2FE", x"C00E84", x"C03A14", x"C065AE", x"C09152", x"C0BD00",
x"C0E8B7", x"C11478", x"C14043", x"C16C18", x"C197F6", x"C1C3DE", x"C1EFCF", x"C21BCA", x"C247CE", x"C273DC",
x"C29FF4", x"C2CC15", x"C2F83F", x"C32473", x"C350B0", x"C37CF7", x"C3A947", x"C3D5A0", x"C40202", x"C42E6E",
x"C45AE3", x"C48761", x"C4B3E8", x"C4E079", x"C50D12", x"C539B5", x"C56661", x"C59315", x"C5BFD3", x"C5EC9A",
x"C6196A", x"C64642", x"C67324", x"C6A00E", x"C6CD01", x"C6F9FD", x"C72702", x"C75410", x"C78126", x"C7AE45",
x"C7DB6D", x"C8089E", x"C835D7", x"C86318", x"C89063", x"C8BDB5", x"C8EB11", x"C91875", x"C945E1", x"C97356",
x"C9A0D3", x"C9CE58", x"C9FBE6", x"CA297C", x"CA571B", x"CA84C2", x"CAB271", x"CAE028", x"CB0DE7", x"CB3BAF",
x"CB697F", x"CB9756", x"CBC536", x"CBF31E", x"CC210E", x"CC4F06", x"CC7D06", x"CCAB0E", x"CCD91E", x"CD0736",
x"CD3555", x"CD637D", x"CD91AC", x"CDBFE3", x"CDEE22", x"CE1C68", x"CE4AB7", x"CE790C", x"CEA76A", x"CED5CF",
x"CF043C", x"CF32B0", x"CF612C", x"CF8FAF", x"CFBE39", x"CFECCC", x"D01B65", x"D04A06", x"D078AE", x"D0A75E",
x"D0D615", x"D104D3", x"D13399", x"D16265", x"D19139", x"D1C014", x"D1EEF6", x"D21DE0", x"D24CD0", x"D27BC7",
x"D2AAC6", x"D2D9CB", x"D308D8", x"D337EB", x"D36705", x"D39626", x"D3C54E", x"D3F47D", x"D423B2", x"D452EF",
x"D48232", x"D4B17B", x"D4E0CC", x"D51023", x"D53F81", x"D56EE5", x"D59E50", x"D5CDC1", x"D5FD39", x"D62CB7",
x"D65C3C", x"D68BC8", x"D6BB59", x"D6EAF1", x"D71A90", x"D74A34", x"D779DF", x"D7A990", x"D7D948", x"D80905",
x"D838C9", x"D86893", x"D89863", x"D8C839", x"D8F815", x"D927F7", x"D957DF", x"D987CD", x"D9B7C1", x"D9E7BB",
x"DA17BB", x"DA47C1", x"DA77CC", x"DAA7DD", x"DAD7F4", x"DB0811", x"DB3834", x"DB685C", x"DB9889", x"DBC8BD",
x"DBF8F6", x"DC2934", x"DC5978", x"DC89C2", x"DCBA11", x"DCEA65", x"DD1ABF", x"DD4B1E", x"DD7B83", x"DDABED",
x"DDDC5C", x"DE0CD0", x"DE3D4A", x"DE6DC9", x"DE9E4D", x"DECED6", x"DEFF65", x"DF2FF8", x"DF6091", x"DF912E",
x"DFC1D1", x"DFF278", x"E02325", x"E053D6", x"E0848C", x"E0B547", x"E0E607", x"E116CC", x"E14795", x"E17864",
x"E1A937", x"E1DA0E", x"E20AEA", x"E23BCB", x"E26CB1", x"E29D9B", x"E2CE89", x"E2FF7C", x"E33074", x"E36170",
x"E39270", x"E3C375", x"E3F47E", x"E4258C", x"E4569E", x"E487B4", x"E4B8CE", x"E4E9EC", x"E51B0F", x"E54C36",
x"E57D61", x"E5AE90", x"E5DFC3", x"E610FA", x"E64235", x"E67374", x"E6A4B7", x"E6D5FE", x"E70748", x"E73897",
x"E769EA", x"E79B40", x"E7CC9A", x"E7FDF8", x"E82F59", x"E860BE", x"E89227", x"E8C393", x"E8F503", x"E92677",
x"E957EE", x"E98968", x"E9BAE6", x"E9EC68", x"EA1DEC", x"EA4F75", x"EA8100", x"EAB28F", x"EAE421", x"EB15B7",
x"EB474F", x"EB78EB", x"EBAA8A", x"EBDC2C", x"EC0DD1", x"EC3F7A", x"EC7125", x"ECA2D3", x"ECD485", x"ED0639",
x"ED37F0", x"ED69AA", x"ED9B67", x"EDCD27", x"EDFEEA", x"EE30AF", x"EE6277", x"EE9442", x"EEC610", x"EEF7E0",
x"EF29B3", x"EF5B88", x"EF8D60", x"EFBF3B", x"EFF118", x"F022F7", x"F054D9", x"F086BE", x"F0B8A5", x"F0EA8E",
x"F11C79", x"F14E67", x"F18057", x"F1B249", x"F1E43E", x"F21634", x"F2482D", x"F27A28", x"F2AC25", x"F2DE24",
x"F31025", x"F34228", x"F3742D", x"F3A634", x"F3D83D", x"F40A48", x"F43C54", x"F46E63", x"F4A073", x"F4D285",
x"F50499", x"F536AE", x"F568C5", x"F59ADE", x"F5CCF8", x"F5FF14", x"F63131", x"F66350", x"F69570", x"F6C792",
x"F6F9B5", x"F72BDA", x"F75E00", x"F79027", x"F7C250", x"F7F47A", x"F826A5", x"F858D1", x"F88AFF", x"F8BD2D",
x"F8EF5D", x"F9218E", x"F953C0", x"F985F3", x"F9B827", x"F9EA5C", x"FA1C92", x"FA4EC9", x"FA8100", x"FAB339",
x"FAE572", x"FB17AC", x"FB49E7", x"FB7C23", x"FBAE5F", x"FBE09C", x"FC12DA", x"FC4518", x"FC7757", x"FCA996",
x"FCDBD6", x"FD0E16", x"FD4057", x"FD7298", x"FDA4DA", x"FDD71C", x"FE095E", x"FE3BA1", x"FE6DE3", x"FEA026",
x"FED26A", x"FF04AD", x"FF36F1", x"FF6935", x"FF9B79", x"FFCDBD",
    -- Pega aquí los 4096 valores desde "seno_lut_4096_q1_23.txt"
    others => (others => '0')
  );

  signal index           : unsigned(27 downto 0) := (others => '0');
  signal offset          : unsigned(11 downto 0);
  signal salida          : signed(23 downto 0);
  signal cuenta_efectiva : unsigned(27 downto 0);
begin

  process(clk)
  begin
    if rising_edge(clk) then
      if new_freq = '1' then
        index <= (others => '0');
      elsif tick = '1' then
        cuenta_efectiva <= shift_left(resize(cuenta_max, 28), 8); -- *256
        index <= index + cuenta_efectiva;
        case index(27 downto 26) is
          when "00" => offset <= index(25 downto 14); salida <= seno_lut(to_integer(offset));
          when "01" => offset <= not index(25 downto 14); salida <= seno_lut(to_integer(offset));
          when "10" => offset <= index(25 downto 14); salida <= -seno_lut(to_integer(offset));
          when others => offset <= not index(25 downto 14); salida <= -seno_lut(to_integer(offset));
        end case;
      end if;
    end if;
  end process;

  gen_seno_out <= std_logic_vector(salida);
end Behavioral;
